module add_round_key(in_matrix, key, out_matrix);
	input [127:0]in_matrix,key;
	output [127:0]out_matrix;
	assign out_matrix = key ^ out_matrix;
endmodule 